-- see Sync.sv handleDidSaveNotification to see how error messages are handled
